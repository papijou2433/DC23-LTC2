* Extracted by KLayout with GF180MCU LVS runset on : 08/11/2023 02:19

.SUBCKT amp Vout1 CLK Vdd Vin2 Vin1 GND
M$1 \$16 Vout1 Vdd Vdd pfet_03v3 L=0.28U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2 \$9 Vin2 \$16 Vdd pfet_03v3 L=0.28U W=10U AS=2.92P AD=3.38P PS=12.92U
+ PD=15.38U
M$7 \$9 \$3 GND GND nfet_03v3 L=0.28U W=7U AS=2.03P AD=1.82P PS=12.06U PD=10.64U
M$14 GND Vout1 \$9 GND nfet_03v3 L=0.28U W=2U AS=0.52P AD=0.7P PS=3.04U PD=4.4U
M$16 \$3 CLK Vdd Vdd pfet_03v3 L=0.28U W=4U AS=1.82P AD=1.82P PS=7.82U PD=7.82U
M$18 \$3 CLK GND GND nfet_03v3 L=0.28U W=4U AS=1.39P AD=1.39P PS=7.78U PD=7.78U
M$22 \$I44 Vin1 Vout1 Vdd pfet_03v3 L=0.28U W=10U AS=3.38P AD=2.92P PS=15.38U
+ PD=12.92U
M$27 Vdd \$9 \$I44 Vdd pfet_03v3 L=0.28U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$28 GND \$9 Vout1 GND nfet_03v3 L=0.28U W=2U AS=0.7P AD=0.52P PS=4.4U PD=3.04U
M$30 GND \$3 Vout1 GND nfet_03v3 L=0.28U W=7U AS=1.82P AD=2.03P PS=10.64U
+ PD=12.06U
.ENDS amp
